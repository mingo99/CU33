typedef logic [`OFM_WIDTH-1:0] sum_t;
typedef logic signed [7:0] mult_t;

typedef logic signed [`OFM_WIDTH-1:0] sum_q[$];
