`include "param.svh"
`include "typedef.svh"
